module div (
		input  wire [7:0] numer,    //  lpm_divide_input.numer
		input  wire [7:0] denom,    //                  .denom
		output wire [7:0] quotient, // lpm_divide_output.quotient
		output wire [7:0] remain    //                  .remain
	);
endmodule

